library verilog;
use verilog.vl_types.all;
entity Data_Memory is
    port(
        rst             : in     vl_logic;
        clk             : in     vl_logic;
        WE              : in     vl_logic;
        A               : in     vl_logic_vector(31 downto 0);
        WD              : in     vl_logic_vector(31 downto 0);
        RD              : out    vl_logic_vector(31 downto 0)
    );
end Data_Memory;
