library verilog;
use verilog.vl_types.all;
entity Test_Bench is
end Test_Bench;
